// soc.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc (
		output wire         bus_clk_clk,                     //              bus_clk.clk
		input  wire [31:0]  ctrl_reg_in_port,                //             ctrl_reg.in_port
		output wire [31:0]  ctrl_reg_out_port,               //                     .out_port
		output wire [31:0]  dma_adr_export,                  //              dma_adr.export
		output wire [31:0]  dma_buf_size_export,             //         dma_buf_size.export
		input  wire [31:0]  dma_status_export,               //           dma_status.export
		input  wire [31:0]  encoder_cnt_export,              //          encoder_cnt.export
		output wire         hps_io_hps_io_emac1_inst_TX_CLK, //               hps_io.hps_io_emac1_inst_TX_CLK
		output wire         hps_io_hps_io_emac1_inst_TXD0,   //                     .hps_io_emac1_inst_TXD0
		output wire         hps_io_hps_io_emac1_inst_TXD1,   //                     .hps_io_emac1_inst_TXD1
		output wire         hps_io_hps_io_emac1_inst_TXD2,   //                     .hps_io_emac1_inst_TXD2
		output wire         hps_io_hps_io_emac1_inst_TXD3,   //                     .hps_io_emac1_inst_TXD3
		input  wire         hps_io_hps_io_emac1_inst_RXD0,   //                     .hps_io_emac1_inst_RXD0
		inout  wire         hps_io_hps_io_emac1_inst_MDIO,   //                     .hps_io_emac1_inst_MDIO
		output wire         hps_io_hps_io_emac1_inst_MDC,    //                     .hps_io_emac1_inst_MDC
		input  wire         hps_io_hps_io_emac1_inst_RX_CTL, //                     .hps_io_emac1_inst_RX_CTL
		output wire         hps_io_hps_io_emac1_inst_TX_CTL, //                     .hps_io_emac1_inst_TX_CTL
		input  wire         hps_io_hps_io_emac1_inst_RX_CLK, //                     .hps_io_emac1_inst_RX_CLK
		input  wire         hps_io_hps_io_emac1_inst_RXD1,   //                     .hps_io_emac1_inst_RXD1
		input  wire         hps_io_hps_io_emac1_inst_RXD2,   //                     .hps_io_emac1_inst_RXD2
		input  wire         hps_io_hps_io_emac1_inst_RXD3,   //                     .hps_io_emac1_inst_RXD3
		inout  wire         hps_io_hps_io_sdio_inst_CMD,     //                     .hps_io_sdio_inst_CMD
		inout  wire         hps_io_hps_io_sdio_inst_D0,      //                     .hps_io_sdio_inst_D0
		inout  wire         hps_io_hps_io_sdio_inst_D1,      //                     .hps_io_sdio_inst_D1
		output wire         hps_io_hps_io_sdio_inst_CLK,     //                     .hps_io_sdio_inst_CLK
		inout  wire         hps_io_hps_io_sdio_inst_D2,      //                     .hps_io_sdio_inst_D2
		inout  wire         hps_io_hps_io_sdio_inst_D3,      //                     .hps_io_sdio_inst_D3
		inout  wire         hps_io_hps_io_usb1_inst_D0,      //                     .hps_io_usb1_inst_D0
		inout  wire         hps_io_hps_io_usb1_inst_D1,      //                     .hps_io_usb1_inst_D1
		inout  wire         hps_io_hps_io_usb1_inst_D2,      //                     .hps_io_usb1_inst_D2
		inout  wire         hps_io_hps_io_usb1_inst_D3,      //                     .hps_io_usb1_inst_D3
		inout  wire         hps_io_hps_io_usb1_inst_D4,      //                     .hps_io_usb1_inst_D4
		inout  wire         hps_io_hps_io_usb1_inst_D5,      //                     .hps_io_usb1_inst_D5
		inout  wire         hps_io_hps_io_usb1_inst_D6,      //                     .hps_io_usb1_inst_D6
		inout  wire         hps_io_hps_io_usb1_inst_D7,      //                     .hps_io_usb1_inst_D7
		input  wire         hps_io_hps_io_usb1_inst_CLK,     //                     .hps_io_usb1_inst_CLK
		output wire         hps_io_hps_io_usb1_inst_STP,     //                     .hps_io_usb1_inst_STP
		input  wire         hps_io_hps_io_usb1_inst_DIR,     //                     .hps_io_usb1_inst_DIR
		input  wire         hps_io_hps_io_usb1_inst_NXT,     //                     .hps_io_usb1_inst_NXT
		output wire         hps_io_hps_io_spim1_inst_CLK,    //                     .hps_io_spim1_inst_CLK
		output wire         hps_io_hps_io_spim1_inst_MOSI,   //                     .hps_io_spim1_inst_MOSI
		input  wire         hps_io_hps_io_spim1_inst_MISO,   //                     .hps_io_spim1_inst_MISO
		output wire         hps_io_hps_io_spim1_inst_SS0,    //                     .hps_io_spim1_inst_SS0
		input  wire         hps_io_hps_io_uart0_inst_RX,     //                     .hps_io_uart0_inst_RX
		output wire         hps_io_hps_io_uart0_inst_TX,     //                     .hps_io_uart0_inst_TX
		inout  wire         hps_io_hps_io_i2c0_inst_SDA,     //                     .hps_io_i2c0_inst_SDA
		inout  wire         hps_io_hps_io_i2c0_inst_SCL,     //                     .hps_io_i2c0_inst_SCL
		inout  wire         hps_io_hps_io_i2c1_inst_SDA,     //                     .hps_io_i2c1_inst_SDA
		inout  wire         hps_io_hps_io_i2c1_inst_SCL,     //                     .hps_io_i2c1_inst_SCL
		inout  wire         hps_io_hps_io_gpio_inst_GPIO09,  //                     .hps_io_gpio_inst_GPIO09
		inout  wire         hps_io_hps_io_gpio_inst_GPIO35,  //                     .hps_io_gpio_inst_GPIO35
		inout  wire         hps_io_hps_io_gpio_inst_GPIO40,  //                     .hps_io_gpio_inst_GPIO40
		inout  wire         hps_io_hps_io_gpio_inst_GPIO53,  //                     .hps_io_gpio_inst_GPIO53
		inout  wire         hps_io_hps_io_gpio_inst_GPIO54,  //                     .hps_io_gpio_inst_GPIO54
		inout  wire         hps_io_hps_io_gpio_inst_GPIO61,  //                     .hps_io_gpio_inst_GPIO61
		input  wire         i_pll_0_refclk_50mhz_clk,        // i_pll_0_refclk_50mhz.clk
		input  wire [31:0]  irq0_irq,                        //                 irq0.irq
		output wire [31:0]  led_clk_on_blue_export,          //      led_clk_on_blue.export
		output wire [31:0]  led_clk_on_green_export,         //     led_clk_on_green.export
		output wire [31:0]  led_clk_on_red_export,           //       led_clk_on_red.export
		output wire [31:0]  lines_cnt_encoder_export,        //    lines_cnt_encoder.export
		output wire [31:0]  lines_delay_export,              //          lines_delay.export
		output wire [14:0]  memory_mem_a,                    //               memory.mem_a
		output wire [2:0]   memory_mem_ba,                   //                     .mem_ba
		output wire         memory_mem_ck,                   //                     .mem_ck
		output wire         memory_mem_ck_n,                 //                     .mem_ck_n
		output wire         memory_mem_cke,                  //                     .mem_cke
		output wire         memory_mem_cs_n,                 //                     .mem_cs_n
		output wire         memory_mem_ras_n,                //                     .mem_ras_n
		output wire         memory_mem_cas_n,                //                     .mem_cas_n
		output wire         memory_mem_we_n,                 //                     .mem_we_n
		output wire         memory_mem_reset_n,              //                     .mem_reset_n
		inout  wire [31:0]  memory_mem_dq,                   //                     .mem_dq
		inout  wire [3:0]   memory_mem_dqs,                  //                     .mem_dqs
		inout  wire [3:0]   memory_mem_dqs_n,                //                     .mem_dqs_n
		output wire         memory_mem_odt,                  //                     .mem_odt
		output wire [3:0]   memory_mem_dm,                   //                     .mem_dm
		input  wire         memory_oct_rzqin,                //                     .oct_rzqin
		output wire         outclk_0_clk,                    //             outclk_0.clk
		output wire         outclk_1_clk,                    //             outclk_1.clk
		input  wire [27:0]  sdram0_address,                  //               sdram0.address
		input  wire [7:0]   sdram0_burstcount,               //                     .burstcount
		output wire         sdram0_waitrequest,              //                     .waitrequest
		output wire [127:0] sdram0_readdata,                 //                     .readdata
		output wire         sdram0_readdatavalid,            //                     .readdatavalid
		input  wire         sdram0_read,                     //                     .read
		input  wire [127:0] sdram0_writedata,                //                     .writedata
		input  wire [15:0]  sdram0_byteenable,               //                     .byteenable
		input  wire         sdram0_write,                    //                     .write
		input  wire [31:0]  status_reg_export,               //           status_reg.export
		input  wire [31:0]  timer_cnt_export                 //            timer_cnt.export
	);

	wire         hps_0_h2f_reset_reset;                                 // hps_0:h2f_rst_n -> [pll_0:rst, rst_controller:reset_in0]
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                       // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                         // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                         // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                        // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                        // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                         // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                           // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                       // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                        // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                        // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                        // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                        // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                         // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                       // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                       // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                          // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                        // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                        // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                        // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                       // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                       // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                       // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                        // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                        // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                         // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                          // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                        // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                        // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                       // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                        // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire         mm_interconnect_0_pio_dma_buf_size_s1_chipselect;      // mm_interconnect_0:pio_dma_buf_size_s1_chipselect -> pio_dma_buf_size:chipselect
	wire  [31:0] mm_interconnect_0_pio_dma_buf_size_s1_readdata;        // pio_dma_buf_size:readdata -> mm_interconnect_0:pio_dma_buf_size_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_dma_buf_size_s1_address;         // mm_interconnect_0:pio_dma_buf_size_s1_address -> pio_dma_buf_size:address
	wire         mm_interconnect_0_pio_dma_buf_size_s1_write;           // mm_interconnect_0:pio_dma_buf_size_s1_write -> pio_dma_buf_size:write_n
	wire  [31:0] mm_interconnect_0_pio_dma_buf_size_s1_writedata;       // mm_interconnect_0:pio_dma_buf_size_s1_writedata -> pio_dma_buf_size:writedata
	wire         mm_interconnect_0_pio_dma_adr_s1_chipselect;           // mm_interconnect_0:pio_dma_adr_s1_chipselect -> pio_dma_adr:chipselect
	wire  [31:0] mm_interconnect_0_pio_dma_adr_s1_readdata;             // pio_dma_adr:readdata -> mm_interconnect_0:pio_dma_adr_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_dma_adr_s1_address;              // mm_interconnect_0:pio_dma_adr_s1_address -> pio_dma_adr:address
	wire         mm_interconnect_0_pio_dma_adr_s1_write;                // mm_interconnect_0:pio_dma_adr_s1_write -> pio_dma_adr:write_n
	wire  [31:0] mm_interconnect_0_pio_dma_adr_s1_writedata;            // mm_interconnect_0:pio_dma_adr_s1_writedata -> pio_dma_adr:writedata
	wire  [31:0] mm_interconnect_0_pio_dma_status_s1_readdata;          // pio_dma_status:readdata -> mm_interconnect_0:pio_dma_status_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_dma_status_s1_address;           // mm_interconnect_0:pio_dma_status_s1_address -> pio_dma_status:address
	wire         mm_interconnect_0_pio_ctrl_reg_s1_chipselect;          // mm_interconnect_0:pio_ctrl_reg_s1_chipselect -> pio_ctrl_reg:chipselect
	wire  [31:0] mm_interconnect_0_pio_ctrl_reg_s1_readdata;            // pio_ctrl_reg:readdata -> mm_interconnect_0:pio_ctrl_reg_s1_readdata
	wire   [2:0] mm_interconnect_0_pio_ctrl_reg_s1_address;             // mm_interconnect_0:pio_ctrl_reg_s1_address -> pio_ctrl_reg:address
	wire         mm_interconnect_0_pio_ctrl_reg_s1_write;               // mm_interconnect_0:pio_ctrl_reg_s1_write -> pio_ctrl_reg:write_n
	wire  [31:0] mm_interconnect_0_pio_ctrl_reg_s1_writedata;           // mm_interconnect_0:pio_ctrl_reg_s1_writedata -> pio_ctrl_reg:writedata
	wire  [31:0] mm_interconnect_0_pio_status_reg_s1_readdata;          // pio_status_reg:readdata -> mm_interconnect_0:pio_status_reg_s1_readdata
	wire   [2:0] mm_interconnect_0_pio_status_reg_s1_address;           // mm_interconnect_0:pio_status_reg_s1_address -> pio_status_reg:address
	wire         mm_interconnect_0_pio_led_clk_on_0_s1_chipselect;      // mm_interconnect_0:pio_led_clk_on_0_s1_chipselect -> pio_led_clk_on_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_clk_on_0_s1_readdata;        // pio_led_clk_on_0:readdata -> mm_interconnect_0:pio_led_clk_on_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_led_clk_on_0_s1_address;         // mm_interconnect_0:pio_led_clk_on_0_s1_address -> pio_led_clk_on_0:address
	wire         mm_interconnect_0_pio_led_clk_on_0_s1_write;           // mm_interconnect_0:pio_led_clk_on_0_s1_write -> pio_led_clk_on_0:write_n
	wire  [31:0] mm_interconnect_0_pio_led_clk_on_0_s1_writedata;       // mm_interconnect_0:pio_led_clk_on_0_s1_writedata -> pio_led_clk_on_0:writedata
	wire         mm_interconnect_0_pio_led_clk_on_1_s1_chipselect;      // mm_interconnect_0:pio_led_clk_on_1_s1_chipselect -> pio_led_clk_on_1:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_clk_on_1_s1_readdata;        // pio_led_clk_on_1:readdata -> mm_interconnect_0:pio_led_clk_on_1_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_led_clk_on_1_s1_address;         // mm_interconnect_0:pio_led_clk_on_1_s1_address -> pio_led_clk_on_1:address
	wire         mm_interconnect_0_pio_led_clk_on_1_s1_write;           // mm_interconnect_0:pio_led_clk_on_1_s1_write -> pio_led_clk_on_1:write_n
	wire  [31:0] mm_interconnect_0_pio_led_clk_on_1_s1_writedata;       // mm_interconnect_0:pio_led_clk_on_1_s1_writedata -> pio_led_clk_on_1:writedata
	wire         mm_interconnect_0_pio_led_clk_on_2_s1_chipselect;      // mm_interconnect_0:pio_led_clk_on_2_s1_chipselect -> pio_led_clk_on_2:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_clk_on_2_s1_readdata;        // pio_led_clk_on_2:readdata -> mm_interconnect_0:pio_led_clk_on_2_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_led_clk_on_2_s1_address;         // mm_interconnect_0:pio_led_clk_on_2_s1_address -> pio_led_clk_on_2:address
	wire         mm_interconnect_0_pio_led_clk_on_2_s1_write;           // mm_interconnect_0:pio_led_clk_on_2_s1_write -> pio_led_clk_on_2:write_n
	wire  [31:0] mm_interconnect_0_pio_led_clk_on_2_s1_writedata;       // mm_interconnect_0:pio_led_clk_on_2_s1_writedata -> pio_led_clk_on_2:writedata
	wire  [31:0] mm_interconnect_0_pio_timer_s1_readdata;               // pio_timer:readdata -> mm_interconnect_0:pio_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_pio_timer_s1_address;                // mm_interconnect_0:pio_timer_s1_address -> pio_timer:address
	wire         mm_interconnect_0_pio_lines_delay_s1_chipselect;       // mm_interconnect_0:pio_lines_delay_s1_chipselect -> pio_lines_delay:chipselect
	wire  [31:0] mm_interconnect_0_pio_lines_delay_s1_readdata;         // pio_lines_delay:readdata -> mm_interconnect_0:pio_lines_delay_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_lines_delay_s1_address;          // mm_interconnect_0:pio_lines_delay_s1_address -> pio_lines_delay:address
	wire         mm_interconnect_0_pio_lines_delay_s1_write;            // mm_interconnect_0:pio_lines_delay_s1_write -> pio_lines_delay:write_n
	wire  [31:0] mm_interconnect_0_pio_lines_delay_s1_writedata;        // mm_interconnect_0:pio_lines_delay_s1_writedata -> pio_lines_delay:writedata
	wire         mm_interconnect_0_pio_lines_cnt_encoder_s1_chipselect; // mm_interconnect_0:pio_lines_cnt_encoder_s1_chipselect -> pio_lines_cnt_encoder:chipselect
	wire  [31:0] mm_interconnect_0_pio_lines_cnt_encoder_s1_readdata;   // pio_lines_cnt_encoder:readdata -> mm_interconnect_0:pio_lines_cnt_encoder_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_lines_cnt_encoder_s1_address;    // mm_interconnect_0:pio_lines_cnt_encoder_s1_address -> pio_lines_cnt_encoder:address
	wire         mm_interconnect_0_pio_lines_cnt_encoder_s1_write;      // mm_interconnect_0:pio_lines_cnt_encoder_s1_write -> pio_lines_cnt_encoder:write_n
	wire  [31:0] mm_interconnect_0_pio_lines_cnt_encoder_s1_writedata;  // mm_interconnect_0:pio_lines_cnt_encoder_s1_writedata -> pio_lines_cnt_encoder:writedata
	wire  [31:0] mm_interconnect_0_pio_encoder_cnt_s1_readdata;         // pio_encoder_cnt:readdata -> mm_interconnect_0:pio_encoder_cnt_s1_readdata
	wire   [2:0] mm_interconnect_0_pio_encoder_cnt_s1_address;          // mm_interconnect_0:pio_encoder_cnt_s1_address -> pio_encoder_cnt:address
	wire  [31:0] hps_0_f2h_irq1_irq;                                    // irq_mapper:sender_irq -> hps_0:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [mm_interconnect_0:pio_dma_buf_size_reset_reset_bridge_in_reset_reset, pio_ctrl_reg:reset_n, pio_dma_adr:reset_n, pio_dma_buf_size:reset_n, pio_dma_status:reset_n, pio_encoder_cnt:reset_n, pio_led_clk_on_0:reset_n, pio_led_clk_on_1:reset_n, pio_led_clk_on_2:reset_n, pio_lines_cnt_encoder:reset_n, pio_lines_delay:reset_n, pio_status_reg:reset_n, pio_timer:reset_n]

	soc_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.mem_a                    (memory_mem_a),                    //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                   //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                   //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                  //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),              //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                   //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                  //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                   //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK), //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL), //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL), //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK), //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),   //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),     //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),    //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),   //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),   //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),    //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),     //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),     //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),     //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),     //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),     //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),  //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),  //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),  //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),  //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),  //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),  //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.f2h_sdram0_clk           (bus_clk_clk),                     //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (sdram0_address),                  //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (sdram0_burstcount),               //                  .burstcount
		.f2h_sdram0_WAITREQUEST   (sdram0_waitrequest),              //                  .waitrequest
		.f2h_sdram0_READDATA      (sdram0_readdata),                 //                  .readdata
		.f2h_sdram0_READDATAVALID (sdram0_readdatavalid),            //                  .readdatavalid
		.f2h_sdram0_READ          (sdram0_read),                     //                  .read
		.f2h_sdram0_WRITEDATA     (sdram0_writedata),                //                  .writedata
		.f2h_sdram0_BYTEENABLE    (sdram0_byteenable),               //                  .byteenable
		.f2h_sdram0_WRITE         (sdram0_write),                    //                  .write
		.h2f_lw_axi_clk           (bus_clk_clk),                     //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0               (irq0_irq),                        //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	soc_pio_ctrl_reg pio_ctrl_reg (
		.clk        (bus_clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_pio_ctrl_reg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_ctrl_reg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_ctrl_reg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_ctrl_reg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_ctrl_reg_s1_readdata),   //                    .readdata
		.in_port    (ctrl_reg_in_port),                             // external_connection.export
		.out_port   (ctrl_reg_out_port)                             //                    .export
	);

	soc_pio_dma_adr pio_dma_adr (
		.clk        (bus_clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pio_dma_adr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_dma_adr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_dma_adr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_dma_adr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_dma_adr_s1_readdata),   //                    .readdata
		.out_port   (dma_adr_export)                               // external_connection.export
	);

	soc_pio_dma_adr pio_dma_buf_size (
		.clk        (bus_clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_pio_dma_buf_size_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_dma_buf_size_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_dma_buf_size_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_dma_buf_size_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_dma_buf_size_s1_readdata),   //                    .readdata
		.out_port   (dma_buf_size_export)                               // external_connection.export
	);

	soc_pio_dma_status pio_dma_status (
		.clk      (bus_clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_pio_dma_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_dma_status_s1_readdata), //                    .readdata
		.in_port  (dma_status_export)                             // external_connection.export
	);

	soc_pio_encoder_cnt pio_encoder_cnt (
		.clk      (bus_clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_pio_encoder_cnt_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_encoder_cnt_s1_readdata), //                    .readdata
		.in_port  (encoder_cnt_export)                             // external_connection.export
	);

	soc_pio_dma_adr pio_led_clk_on_0 (
		.clk        (bus_clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_clk_on_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_clk_on_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_clk_on_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_clk_on_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_clk_on_0_s1_readdata),   //                    .readdata
		.out_port   (led_clk_on_red_export)                             // external_connection.export
	);

	soc_pio_dma_adr pio_led_clk_on_1 (
		.clk        (bus_clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_clk_on_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_clk_on_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_clk_on_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_clk_on_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_clk_on_1_s1_readdata),   //                    .readdata
		.out_port   (led_clk_on_green_export)                           // external_connection.export
	);

	soc_pio_dma_adr pio_led_clk_on_2 (
		.clk        (bus_clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_clk_on_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_clk_on_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_clk_on_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_clk_on_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_clk_on_2_s1_readdata),   //                    .readdata
		.out_port   (led_clk_on_blue_export)                            // external_connection.export
	);

	soc_pio_dma_adr pio_lines_cnt_encoder (
		.clk        (bus_clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (mm_interconnect_0_pio_lines_cnt_encoder_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_lines_cnt_encoder_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_lines_cnt_encoder_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_lines_cnt_encoder_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_lines_cnt_encoder_s1_readdata),   //                    .readdata
		.out_port   (lines_cnt_encoder_export)                               // external_connection.export
	);

	soc_pio_dma_adr pio_lines_delay (
		.clk        (bus_clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_pio_lines_delay_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_lines_delay_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_lines_delay_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_lines_delay_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_lines_delay_s1_readdata),   //                    .readdata
		.out_port   (lines_delay_export)                               // external_connection.export
	);

	soc_pio_encoder_cnt pio_status_reg (
		.clk      (bus_clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_pio_status_reg_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_status_reg_s1_readdata), //                    .readdata
		.in_port  (status_reg_export)                             // external_connection.export
	);

	soc_pio_encoder_cnt pio_timer (
		.clk      (bus_clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_pio_timer_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_timer_s1_readdata), //                    .readdata
		.in_port  (timer_cnt_export)                         // external_connection.export
	);

	soc_pll_0 pll_0 (
		.refclk   (i_pll_0_refclk_50mhz_clk), //  refclk.clk
		.rst      (~hps_0_h2f_reset_reset),   //   reset.reset
		.outclk_0 (bus_clk_clk),              // outclk0.clk
		.outclk_1 (outclk_0_clk),             // outclk1.clk
		.outclk_2 (outclk_1_clk),             // outclk2.clk
		.locked   ()                          // (terminated)
	);

	soc_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                       (hps_0_h2f_lw_axi_master_awid),                          //                      hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                     (hps_0_h2f_lw_axi_master_awaddr),                        //                                             .awaddr
		.hps_0_h2f_lw_axi_master_awlen                      (hps_0_h2f_lw_axi_master_awlen),                         //                                             .awlen
		.hps_0_h2f_lw_axi_master_awsize                     (hps_0_h2f_lw_axi_master_awsize),                        //                                             .awsize
		.hps_0_h2f_lw_axi_master_awburst                    (hps_0_h2f_lw_axi_master_awburst),                       //                                             .awburst
		.hps_0_h2f_lw_axi_master_awlock                     (hps_0_h2f_lw_axi_master_awlock),                        //                                             .awlock
		.hps_0_h2f_lw_axi_master_awcache                    (hps_0_h2f_lw_axi_master_awcache),                       //                                             .awcache
		.hps_0_h2f_lw_axi_master_awprot                     (hps_0_h2f_lw_axi_master_awprot),                        //                                             .awprot
		.hps_0_h2f_lw_axi_master_awvalid                    (hps_0_h2f_lw_axi_master_awvalid),                       //                                             .awvalid
		.hps_0_h2f_lw_axi_master_awready                    (hps_0_h2f_lw_axi_master_awready),                       //                                             .awready
		.hps_0_h2f_lw_axi_master_wid                        (hps_0_h2f_lw_axi_master_wid),                           //                                             .wid
		.hps_0_h2f_lw_axi_master_wdata                      (hps_0_h2f_lw_axi_master_wdata),                         //                                             .wdata
		.hps_0_h2f_lw_axi_master_wstrb                      (hps_0_h2f_lw_axi_master_wstrb),                         //                                             .wstrb
		.hps_0_h2f_lw_axi_master_wlast                      (hps_0_h2f_lw_axi_master_wlast),                         //                                             .wlast
		.hps_0_h2f_lw_axi_master_wvalid                     (hps_0_h2f_lw_axi_master_wvalid),                        //                                             .wvalid
		.hps_0_h2f_lw_axi_master_wready                     (hps_0_h2f_lw_axi_master_wready),                        //                                             .wready
		.hps_0_h2f_lw_axi_master_bid                        (hps_0_h2f_lw_axi_master_bid),                           //                                             .bid
		.hps_0_h2f_lw_axi_master_bresp                      (hps_0_h2f_lw_axi_master_bresp),                         //                                             .bresp
		.hps_0_h2f_lw_axi_master_bvalid                     (hps_0_h2f_lw_axi_master_bvalid),                        //                                             .bvalid
		.hps_0_h2f_lw_axi_master_bready                     (hps_0_h2f_lw_axi_master_bready),                        //                                             .bready
		.hps_0_h2f_lw_axi_master_arid                       (hps_0_h2f_lw_axi_master_arid),                          //                                             .arid
		.hps_0_h2f_lw_axi_master_araddr                     (hps_0_h2f_lw_axi_master_araddr),                        //                                             .araddr
		.hps_0_h2f_lw_axi_master_arlen                      (hps_0_h2f_lw_axi_master_arlen),                         //                                             .arlen
		.hps_0_h2f_lw_axi_master_arsize                     (hps_0_h2f_lw_axi_master_arsize),                        //                                             .arsize
		.hps_0_h2f_lw_axi_master_arburst                    (hps_0_h2f_lw_axi_master_arburst),                       //                                             .arburst
		.hps_0_h2f_lw_axi_master_arlock                     (hps_0_h2f_lw_axi_master_arlock),                        //                                             .arlock
		.hps_0_h2f_lw_axi_master_arcache                    (hps_0_h2f_lw_axi_master_arcache),                       //                                             .arcache
		.hps_0_h2f_lw_axi_master_arprot                     (hps_0_h2f_lw_axi_master_arprot),                        //                                             .arprot
		.hps_0_h2f_lw_axi_master_arvalid                    (hps_0_h2f_lw_axi_master_arvalid),                       //                                             .arvalid
		.hps_0_h2f_lw_axi_master_arready                    (hps_0_h2f_lw_axi_master_arready),                       //                                             .arready
		.hps_0_h2f_lw_axi_master_rid                        (hps_0_h2f_lw_axi_master_rid),                           //                                             .rid
		.hps_0_h2f_lw_axi_master_rdata                      (hps_0_h2f_lw_axi_master_rdata),                         //                                             .rdata
		.hps_0_h2f_lw_axi_master_rresp                      (hps_0_h2f_lw_axi_master_rresp),                         //                                             .rresp
		.hps_0_h2f_lw_axi_master_rlast                      (hps_0_h2f_lw_axi_master_rlast),                         //                                             .rlast
		.hps_0_h2f_lw_axi_master_rvalid                     (hps_0_h2f_lw_axi_master_rvalid),                        //                                             .rvalid
		.hps_0_h2f_lw_axi_master_rready                     (hps_0_h2f_lw_axi_master_rready),                        //                                             .rready
		.pll_0_outclk0_clk                                  (bus_clk_clk),                                           //                                pll_0_outclk0.clk
		.pio_dma_buf_size_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // pio_dma_buf_size_reset_reset_bridge_in_reset.reset
		.pio_ctrl_reg_s1_address                            (mm_interconnect_0_pio_ctrl_reg_s1_address),             //                              pio_ctrl_reg_s1.address
		.pio_ctrl_reg_s1_write                              (mm_interconnect_0_pio_ctrl_reg_s1_write),               //                                             .write
		.pio_ctrl_reg_s1_readdata                           (mm_interconnect_0_pio_ctrl_reg_s1_readdata),            //                                             .readdata
		.pio_ctrl_reg_s1_writedata                          (mm_interconnect_0_pio_ctrl_reg_s1_writedata),           //                                             .writedata
		.pio_ctrl_reg_s1_chipselect                         (mm_interconnect_0_pio_ctrl_reg_s1_chipselect),          //                                             .chipselect
		.pio_dma_adr_s1_address                             (mm_interconnect_0_pio_dma_adr_s1_address),              //                               pio_dma_adr_s1.address
		.pio_dma_adr_s1_write                               (mm_interconnect_0_pio_dma_adr_s1_write),                //                                             .write
		.pio_dma_adr_s1_readdata                            (mm_interconnect_0_pio_dma_adr_s1_readdata),             //                                             .readdata
		.pio_dma_adr_s1_writedata                           (mm_interconnect_0_pio_dma_adr_s1_writedata),            //                                             .writedata
		.pio_dma_adr_s1_chipselect                          (mm_interconnect_0_pio_dma_adr_s1_chipselect),           //                                             .chipselect
		.pio_dma_buf_size_s1_address                        (mm_interconnect_0_pio_dma_buf_size_s1_address),         //                          pio_dma_buf_size_s1.address
		.pio_dma_buf_size_s1_write                          (mm_interconnect_0_pio_dma_buf_size_s1_write),           //                                             .write
		.pio_dma_buf_size_s1_readdata                       (mm_interconnect_0_pio_dma_buf_size_s1_readdata),        //                                             .readdata
		.pio_dma_buf_size_s1_writedata                      (mm_interconnect_0_pio_dma_buf_size_s1_writedata),       //                                             .writedata
		.pio_dma_buf_size_s1_chipselect                     (mm_interconnect_0_pio_dma_buf_size_s1_chipselect),      //                                             .chipselect
		.pio_dma_status_s1_address                          (mm_interconnect_0_pio_dma_status_s1_address),           //                            pio_dma_status_s1.address
		.pio_dma_status_s1_readdata                         (mm_interconnect_0_pio_dma_status_s1_readdata),          //                                             .readdata
		.pio_encoder_cnt_s1_address                         (mm_interconnect_0_pio_encoder_cnt_s1_address),          //                           pio_encoder_cnt_s1.address
		.pio_encoder_cnt_s1_readdata                        (mm_interconnect_0_pio_encoder_cnt_s1_readdata),         //                                             .readdata
		.pio_led_clk_on_0_s1_address                        (mm_interconnect_0_pio_led_clk_on_0_s1_address),         //                          pio_led_clk_on_0_s1.address
		.pio_led_clk_on_0_s1_write                          (mm_interconnect_0_pio_led_clk_on_0_s1_write),           //                                             .write
		.pio_led_clk_on_0_s1_readdata                       (mm_interconnect_0_pio_led_clk_on_0_s1_readdata),        //                                             .readdata
		.pio_led_clk_on_0_s1_writedata                      (mm_interconnect_0_pio_led_clk_on_0_s1_writedata),       //                                             .writedata
		.pio_led_clk_on_0_s1_chipselect                     (mm_interconnect_0_pio_led_clk_on_0_s1_chipselect),      //                                             .chipselect
		.pio_led_clk_on_1_s1_address                        (mm_interconnect_0_pio_led_clk_on_1_s1_address),         //                          pio_led_clk_on_1_s1.address
		.pio_led_clk_on_1_s1_write                          (mm_interconnect_0_pio_led_clk_on_1_s1_write),           //                                             .write
		.pio_led_clk_on_1_s1_readdata                       (mm_interconnect_0_pio_led_clk_on_1_s1_readdata),        //                                             .readdata
		.pio_led_clk_on_1_s1_writedata                      (mm_interconnect_0_pio_led_clk_on_1_s1_writedata),       //                                             .writedata
		.pio_led_clk_on_1_s1_chipselect                     (mm_interconnect_0_pio_led_clk_on_1_s1_chipselect),      //                                             .chipselect
		.pio_led_clk_on_2_s1_address                        (mm_interconnect_0_pio_led_clk_on_2_s1_address),         //                          pio_led_clk_on_2_s1.address
		.pio_led_clk_on_2_s1_write                          (mm_interconnect_0_pio_led_clk_on_2_s1_write),           //                                             .write
		.pio_led_clk_on_2_s1_readdata                       (mm_interconnect_0_pio_led_clk_on_2_s1_readdata),        //                                             .readdata
		.pio_led_clk_on_2_s1_writedata                      (mm_interconnect_0_pio_led_clk_on_2_s1_writedata),       //                                             .writedata
		.pio_led_clk_on_2_s1_chipselect                     (mm_interconnect_0_pio_led_clk_on_2_s1_chipselect),      //                                             .chipselect
		.pio_lines_cnt_encoder_s1_address                   (mm_interconnect_0_pio_lines_cnt_encoder_s1_address),    //                     pio_lines_cnt_encoder_s1.address
		.pio_lines_cnt_encoder_s1_write                     (mm_interconnect_0_pio_lines_cnt_encoder_s1_write),      //                                             .write
		.pio_lines_cnt_encoder_s1_readdata                  (mm_interconnect_0_pio_lines_cnt_encoder_s1_readdata),   //                                             .readdata
		.pio_lines_cnt_encoder_s1_writedata                 (mm_interconnect_0_pio_lines_cnt_encoder_s1_writedata),  //                                             .writedata
		.pio_lines_cnt_encoder_s1_chipselect                (mm_interconnect_0_pio_lines_cnt_encoder_s1_chipselect), //                                             .chipselect
		.pio_lines_delay_s1_address                         (mm_interconnect_0_pio_lines_delay_s1_address),          //                           pio_lines_delay_s1.address
		.pio_lines_delay_s1_write                           (mm_interconnect_0_pio_lines_delay_s1_write),            //                                             .write
		.pio_lines_delay_s1_readdata                        (mm_interconnect_0_pio_lines_delay_s1_readdata),         //                                             .readdata
		.pio_lines_delay_s1_writedata                       (mm_interconnect_0_pio_lines_delay_s1_writedata),        //                                             .writedata
		.pio_lines_delay_s1_chipselect                      (mm_interconnect_0_pio_lines_delay_s1_chipselect),       //                                             .chipselect
		.pio_status_reg_s1_address                          (mm_interconnect_0_pio_status_reg_s1_address),           //                            pio_status_reg_s1.address
		.pio_status_reg_s1_readdata                         (mm_interconnect_0_pio_status_reg_s1_readdata),          //                                             .readdata
		.pio_timer_s1_address                               (mm_interconnect_0_pio_timer_s1_address),                //                                 pio_timer_s1.address
		.pio_timer_s1_readdata                              (mm_interconnect_0_pio_timer_s1_readdata)                //                                             .readdata
	);

	soc_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (bus_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
